`ifndef BPB_VH
`define BPB_VH

`timescale 1ns / 1ps

// number of entries
`define BPB_E 8
// index bits
`define BPB_T 10

`endif